library verilog;
use verilog.vl_types.all;
entity multiplicadorPor9_vlg_vec_tst is
end multiplicadorPor9_vlg_vec_tst;
