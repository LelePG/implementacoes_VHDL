library verilog;
use verilog.vl_types.all;
entity processador_vlg_check_tst is
    port(
        saidaTeste      : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end processador_vlg_check_tst;
