library verilog;
use verilog.vl_types.all;
entity multiplicadorMatricial_vlg_vec_tst is
end multiplicadorMatricial_vlg_vec_tst;
