library verilog;
use verilog.vl_types.all;
entity debug_vlg_vec_tst is
end debug_vlg_vec_tst;
