library verilog;
use verilog.vl_types.all;
entity multiplicadorSequencial_vlg_vec_tst is
end multiplicadorSequencial_vlg_vec_tst;
